
module Adder(input[31:0] a, input[31:0] b, output[31:0] f);
	assign f = a + b;
endmodule